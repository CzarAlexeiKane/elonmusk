conectix             *D}�vbox  Wi2k    @      @  �?   ���d9��a�'C�����#                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������             �    ���}                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                        conectix             *D}�vbox  Wi2k    @      @  �?   ���d9��a�'C�����#                                                                                                                                                                                                                                                                                                                                                                                                                                            